module main

fn main() {
	print_hello_from_lua()
}
